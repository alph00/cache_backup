module mmu(

);

endmodule